library verilog;
use verilog.vl_types.all;
entity choin_vlg_vec_tst is
end choin_vlg_vec_tst;
